
//----------------------------------------------------------------
// Declare
//----------------------------------------------------------------

// Using UTF-8.
// System Verilog
// ALL RIGHTS RESERVED BY ClARK.

module decoder_3to8

//----------------------------------------------------------------
// Ports
//----------------------------------------------------------------

(
     code_i
    ,decode_o
);

    // Inputs
    input logic [2:0] code_i;

    // Outputs
    output logic [7:0] decode_o;

//----------------------------------------------------------------
// Registers / Wires / Params / Includes
//----------------------------------------------------------------

parameter ONE_8B = 8'b0000_0001;

//----------------------------------------------------------------
// Test Bench
//----------------------------------------------------------------

// reg [2:0] code_i = 3'bxxx;
// integer row = 0;

// initial begin
//     for (row = 0; row <= 8; row = row + 1) begin
//         #(10) code_i = row;
//     end
// end

//----------------------------------------------------------------
// Circuits
//----------------------------------------------------------------

always_comb begin
    if (code_i == 0)
        decode_o = '0;
    else if (0 < code_i && code_i <= '1)
        decode_o = ONE_8B << (code_i - 1);
    else
        decode_o = 'x;
end

endmodule
